module video_top
    (
        input [12:0] ADDRESS,
        input IE,
        input [1:0] COLOUR,
        input PALETTE_SW,
        input             I_clk           ,
        input             I_rst           ,
        input             I_key           ,
        output            running         ,
        output            O_tmds_clk_p    ,
        output            O_tmds_clk_n    ,
        output     [2:0]  O_tmds_data_p   ,
        output     [2:0]  O_tmds_data_n   
    );

    wire [12:0] pixel_address;
    wire [1:0] pixel_colour;

    wire [1:0] palette;

    wire [23:0] bgcolour;

    assign      I_rst_n = ~I_rst;

    reg  [1:0]  KEY_sync;

    reg  [31:0] run_cnt;
    wire        running;
    wire        I_rst_n;

    reg [1:0] KEY_sync;
    always @(posedge pix_clk or negedge hdmi4_rst_n) begin
        if (!hdmi4_rst_n)    
            KEY_sync <= 2'b00;
        else                 
            KEY_sync <= {KEY_sync[0], I_key};
    end


    wire KEY_pressed =  KEY_sync[0] & ~KEY_sync[1];

    reg [2:0]   mode_reg;

    always @(posedge pix_clk or negedge hdmi4_rst_n) begin
        if (!hdmi4_rst_n)      
            mode_reg <= 3'd0;
        else if (KEY_pressed)   
            mode_reg <= mode_reg + 3'd1;
        else                   
            mode_reg <= mode_reg;
    end


    //--------------------------
    wire        tp0_vs_in  ;
    wire        tp0_hs_in  ;
    wire        tp0_de_in ;
    wire [ 7:0] tp0_data_r/*synthesis syn_keep=1*/;
    wire [ 7:0] tp0_data_g/*synthesis syn_keep=1*/;
    wire [ 7:0] tp0_data_b/*synthesis syn_keep=1*/;

    reg         vs_r;
    reg  [9:0]  cnt_vs;

    //------------------------------------
    //HDMI4 TX
    wire serial_clk;
    wire pll_lock;

    wire hdmi4_rst_n;

    wire pix_clk;

    always @(posedge I_clk or negedge I_rst_n) //I_clk
    begin
        if(!I_rst_n)
            run_cnt <= 32'd0;
        else if(run_cnt >= 32'd27_000_000)
            run_cnt <= 32'd0;
        else
            run_cnt <= run_cnt + 1'b1;
    end

    assign  running = (run_cnt < 32'd14_000_000) ? 1'b1 : 1'b0;

    testpattern testpattern_inst
    (
        .I_pxl_clk   (pix_clk            ),//pixel clock
        .I_rst_n     (hdmi4_rst_n        ),//low active 
        .I_mode      (mode_reg           ),//data select
        .I_single_r  (8'd0               ),
        .I_single_g  (8'd255             ),
        .I_single_b  (8'd0               ),                  //800x600    //1024x768   //1280x720    
        .I_h_total   (12'd1650           ),//hor total time  // 12'd1056  // 12'd1344  // 12'd1650  
        .I_h_sync    (12'd40             ),//hor sync time   // 12'd128   // 12'd136   // 12'd40    
        .I_h_bporch  (12'd220            ),//hor back porch  // 12'd88    // 12'd160   // 12'd220   
        .I_h_res     (12'd1280           ),//hor resolution  // 12'd800   // 12'd1024  // 12'd1280  
        .I_v_total   (12'd750            ),//ver total time  // 12'd628   // 12'd806   // 12'd750    
        .I_v_sync    (12'd5              ),//ver sync time   // 12'd4     // 12'd6     // 12'd5     
        .I_v_bporch  (12'd20             ),//ver back porch  // 12'd23    // 12'd29    // 12'd20    
        .I_v_res     (12'd720            ),//ver resolution  // 12'd600   // 12'd768   // 12'd720    
        .I_hs_pol    (1'b1               ),//HS polarity , 0:negetive ploarity，1：positive polarity
        .I_vs_pol    (1'b1               ),//VS polarity , 0:negetive ploarity，1：positive polarity
        .O_de        (tp0_de_in          ),   
        .O_hs        (tp0_hs_in          ),
        .O_vs        (tp0_vs_in          ),
        .O_data_r    (tp0_data_r         ),   
        .O_data_g    (tp0_data_g         ),
        .O_data_b    (tp0_data_b         ),
        .pixel_colour(pixel_colour),
        .pixel_address(pixel_address),
        .bgcolour(bgcolour),
        .palette(palette)
    );

    frame_buffer fb (
        .clk(I_clk),
        .address(ADDRESS),
        .addr_internal(pixel_address),
        .colour(COLOUR),
        .IE(IE),
        .dataOut(pixel_colour),
        .bgcolour(bgcolour)
    );

    palette_sw sw1 (
        .palette(palette),
        .sw(PALETTE_SW),
        .clk(I_clk)
    );

    always@(posedge pix_clk) begin
        vs_r<=tp0_vs_in;
    end

    always@(posedge pix_clk or negedge hdmi4_rst_n)
    begin
        if(!hdmi4_rst_n)
            cnt_vs<=0;
        else if(vs_r && !tp0_vs_in) //vKEY4 falling edge
            cnt_vs<=cnt_vs+1'b1;
    end 

    TMDS_rPLL u_tmds_rpll
    (.clkin     (I_clk     )     //input clk 
    ,.clkout    (serial_clk)     //output clk 
    ,.lock      (pll_lock  )     //output lock
    );

    assign hdmi4_rst_n = I_rst_n & pll_lock;

    CLKDIV u_clkdiv
    (.RESETN(hdmi4_rst_n)
    ,.HCLKIN(serial_clk) //clk  x5
    ,.CLKOUT(pix_clk)    //clk  x1
    ,.CALIB (1'b1)
    );
    defparam u_clkdiv.DIV_MODE="5";
    defparam u_clkdiv.GSREN="false";

    DVI_TX_Top DVI_TX_Top_inst
    (
        .I_rst_n       (hdmi4_rst_n   ),  //asynchronous reset, low active
        .I_serial_clk  (serial_clk    ),
        .I_rgb_clk     (pix_clk       ),  //pixel clock
        .I_rgb_vs      (tp0_vs_in     ), 
        .I_rgb_hs      (tp0_hs_in     ),    
        .I_rgb_de      (tp0_de_in     ), 
        .I_rgb_r       (  tp0_data_r ),  //tp0_data_r
        .I_rgb_g       (  tp0_data_g  ),  
        .I_rgb_b       (  tp0_data_b  ),  
        .O_tmds_clk_p  (O_tmds_clk_p  ),
        .O_tmds_clk_n  (O_tmds_clk_n  ),
        .O_tmds_data_p (O_tmds_data_p ),  //{r,g,b}
        .O_tmds_data_n (O_tmds_data_n )
    );

    key_led_ctrl key_led_ctrl_inst
    (
        .I_rst_n       (hdmi4_rst_n   ),
        .I_clk         (pix_clk       ), 
        .I_key         (I_key         )
    );

endmodule